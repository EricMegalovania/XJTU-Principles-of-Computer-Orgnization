`include "defines.v"

// 指令存储器模块
module inst_memory(
    input wire [`ADDR_LEN-1:0] addr,   // 指令地址
    output wire [`INSTR_LEN-1:0] inst  // 读出的指令
);
    
    // 256条指令的指令存储器
    reg [`INSTR_LEN-1:0] inst_mem [0:255];
    
    // 初始化测试指令
    initial begin
        inst_mem[0]  = 32'b001101_00000_00000_0000_0000_0000_0000;
        inst_mem[1]  = 32'b001000_00000_00001_0000_0000_0000_0001;
        inst_mem[2]  = 32'b001101_00000_00010_0000_0000_0000_0010;
        inst_mem[3]  = 32'b000000_00001_00010_00011_00000_100000;
        inst_mem[4]  = 32'b000000_00010_00001_00100_00000_100010;
        inst_mem[5]  = 32'b000100_00011_00100_0000_0000_0000_0100;
        inst_mem[6]  = 32'b000000_00001_00010_00101_00000_100101;
        inst_mem[7]  = 32'b000100_00011_00101_0000_0000_0000_0010;
        inst_mem[8]  = 32'b000010_0000_0000_0000_0000_0000_0000_00;
        inst_mem[9]  = 32'b000010_0000_0000_0000_0000_0000_0010_11;
        inst_mem[10] = 32'b000010_0000_0000_0000_0000_0000_0000_00;
        inst_mem[11] = 32'b000000_00101_00010_00110_00000_100100;
        inst_mem[12] = 32'b000100_00001_00110_0000_0000_0000_0011;
        inst_mem[13] = 32'b000010_0000_0000_0000_0000_0000_0000_00;
        inst_mem[14] = 32'b000010_0000_0000_0000_0000_0000_0000_00;
        inst_mem[15] = 32'b101011_00001_00110_0000_0000_0000_1111;
        inst_mem[16] = 32'b100011_00111_00101_0000_0000_0000_1101;
    end
    
    // 读取指令, 每条指令32位占4字节, 所以地址需要除以4
    assign inst = inst_mem[addr[`ADDR_LEN-1:2]];
    
endmodule
